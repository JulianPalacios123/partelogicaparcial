-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.1.0 Build 162 10/23/2013 SJ Web Edition"
-- CREATED		"Mon Dec 12 00:51:36 2022"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY sietesegmentos IS 
	PORT
	(
		A0 :  IN  STD_LOGIC;
		B0 :  IN  STD_LOGIC;
		C0 :  IN  STD_LOGIC;
		D0 :  IN  STD_LOGIC;
		a :  OUT  STD_LOGIC;
		b :  OUT  STD_LOGIC;
		c :  OUT  STD_LOGIC;
		d :  OUT  STD_LOGIC;
		e :  OUT  STD_LOGIC;
		f :  OUT  STD_LOGIC;
		g :  OUT  STD_LOGIC
	);
END sietesegmentos;

ARCHITECTURE bdf_type OF sietesegmentos IS 

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;


BEGIN 



SYNTHESIZED_WIRE_18 <= SYNTHESIZED_WIRE_0 OR SYNTHESIZED_WIRE_1;


SYNTHESIZED_WIRE_1 <= C0 OR A0;


SYNTHESIZED_WIRE_22 <= NOT(D0);



SYNTHESIZED_WIRE_2 <= C0 AND D0;


SYNTHESIZED_WIRE_17 <= NOT(A0);



SYNTHESIZED_WIRE_30 <= SYNTHESIZED_WIRE_2 OR SYNTHESIZED_WIRE_3 OR SYNTHESIZED_WIRE_4;


SYNTHESIZED_WIRE_37 <= A0 OR SYNTHESIZED_WIRE_5 OR D0 OR B0;


SYNTHESIZED_WIRE_5 <= NOT(C0);



SYNTHESIZED_WIRE_9 <= NOT(B0);



SYNTHESIZED_WIRE_11 <= NOT(B0);



SYNTHESIZED_WIRE_6 <= NOT(C0);



SYNTHESIZED_WIRE_12 <= NOT(D0);



SYNTHESIZED_WIRE_10 <= NOT(D0);



SYNTHESIZED_WIRE_13 <= B0 AND SYNTHESIZED_WIRE_6 AND D0;


SYNTHESIZED_WIRE_39 <= SYNTHESIZED_WIRE_7 AND SYNTHESIZED_WIRE_8;


SYNTHESIZED_WIRE_16 <= SYNTHESIZED_WIRE_9 AND SYNTHESIZED_WIRE_10;


SYNTHESIZED_WIRE_14 <= SYNTHESIZED_WIRE_11 AND C0;


SYNTHESIZED_WIRE_15 <= C0 AND SYNTHESIZED_WIRE_12;


SYNTHESIZED_WIRE_38 <= SYNTHESIZED_WIRE_13 OR SYNTHESIZED_WIRE_14 OR SYNTHESIZED_WIRE_15 OR SYNTHESIZED_WIRE_16;


SYNTHESIZED_WIRE_19 <= SYNTHESIZED_WIRE_17 AND C0;


a <= NOT(SYNTHESIZED_WIRE_18);



SYNTHESIZED_WIRE_8 <= SYNTHESIZED_WIRE_19 OR SYNTHESIZED_WIRE_20;


SYNTHESIZED_WIRE_20 <= SYNTHESIZED_WIRE_21 AND SYNTHESIZED_WIRE_22;


SYNTHESIZED_WIRE_23 <= NOT(C0);



SYNTHESIZED_WIRE_24 <= NOT(D0);



SYNTHESIZED_WIRE_7 <= NOT(D0);



SYNTHESIZED_WIRE_26 <= NOT(D0);



SYNTHESIZED_WIRE_25 <= NOT(C0);



SYNTHESIZED_WIRE_31 <= NOT(B0);



SYNTHESIZED_WIRE_27 <= SYNTHESIZED_WIRE_23 AND SYNTHESIZED_WIRE_24;


SYNTHESIZED_WIRE_29 <= B0 AND SYNTHESIZED_WIRE_25;


SYNTHESIZED_WIRE_28 <= B0 AND SYNTHESIZED_WIRE_26;


SYNTHESIZED_WIRE_40 <= SYNTHESIZED_WIRE_27 OR SYNTHESIZED_WIRE_28 OR A0 OR SYNTHESIZED_WIRE_29;


b <= NOT(SYNTHESIZED_WIRE_30);



SYNTHESIZED_WIRE_36 <= NOT(D0);



SYNTHESIZED_WIRE_32 <= NOT(C0);



SYNTHESIZED_WIRE_0 <= NOT(B0 XOR D0);


SYNTHESIZED_WIRE_33 <= SYNTHESIZED_WIRE_31 AND C0;


SYNTHESIZED_WIRE_35 <= B0 AND SYNTHESIZED_WIRE_32;


SYNTHESIZED_WIRE_41 <= SYNTHESIZED_WIRE_33 OR SYNTHESIZED_WIRE_34 OR A0 OR SYNTHESIZED_WIRE_35;


SYNTHESIZED_WIRE_34 <= C0 AND SYNTHESIZED_WIRE_36;


c <= NOT(SYNTHESIZED_WIRE_37);



d <= NOT(SYNTHESIZED_WIRE_38);



e <= NOT(SYNTHESIZED_WIRE_39);



f <= NOT(SYNTHESIZED_WIRE_40);



g <= NOT(SYNTHESIZED_WIRE_41);



SYNTHESIZED_WIRE_21 <= NOT(B0);



SYNTHESIZED_WIRE_42 <= NOT(C0);



SYNTHESIZED_WIRE_43 <= NOT(D0);



SYNTHESIZED_WIRE_3 <= NOT(B0);



SYNTHESIZED_WIRE_4 <= SYNTHESIZED_WIRE_42 AND SYNTHESIZED_WIRE_43;


END bdf_type;