-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.1.0 Build 162 10/23/2013 SJ Web Edition"
-- CREATED		"Thu Dec 15 16:12:12 2022"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY parcial_digitales IS 
	PORT
	(
		S0 :  IN  STD_LOGIC;
		S1 :  IN  STD_LOGIC;
		A0 :  IN  STD_LOGIC;
		B0 :  IN  STD_LOGIC;
		B1 :  IN  STD_LOGIC;
		A1 :  IN  STD_LOGIC;
		B2 :  IN  STD_LOGIC;
		A2 :  IN  STD_LOGIC;
		A3 :  IN  STD_LOGIC;
		B3 :  IN  STD_LOGIC;
		cin :  IN  STD_LOGIC;
		F0 :  OUT  STD_LOGIC;
		F1 :  OUT  STD_LOGIC;
		F2 :  OUT  STD_LOGIC;
		F3 :  OUT  STD_LOGIC;
		C0 :  OUT  STD_LOGIC;
		b :  OUT  STD_LOGIC;
		c :  OUT  STD_LOGIC;
		d :  OUT  STD_LOGIC;
		e :  OUT  STD_LOGIC;
		f :  OUT  STD_LOGIC;
		g :  OUT  STD_LOGIC;
		a :  OUT  STD_LOGIC
	);
END parcial_digitales;

ARCHITECTURE bdf_type OF parcial_digitales IS 

ATTRIBUTE black_box : BOOLEAN;
ATTRIBUTE noopt : BOOLEAN;

COMPONENT \21mux_10\
	PORT(S : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 A : IN STD_LOGIC;
		 Y : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \21mux_10\: COMPONENT IS true;
ATTRIBUTE noopt OF \21mux_10\: COMPONENT IS true;

COMPONENT \21mux_11\
	PORT(S : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 A : IN STD_LOGIC;
		 Y : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \21mux_11\: COMPONENT IS true;
ATTRIBUTE noopt OF \21mux_11\: COMPONENT IS true;

COMPONENT \21mux_12\
	PORT(S : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 A : IN STD_LOGIC;
		 Y : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \21mux_12\: COMPONENT IS true;
ATTRIBUTE noopt OF \21mux_12\: COMPONENT IS true;

COMPONENT \21mux_13\
	PORT(S : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 A : IN STD_LOGIC;
		 Y : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \21mux_13\: COMPONENT IS true;
ATTRIBUTE noopt OF \21mux_13\: COMPONENT IS true;

COMPONENT \21mux_2\
	PORT(S : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 A : IN STD_LOGIC;
		 Y : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \21mux_2\: COMPONENT IS true;
ATTRIBUTE noopt OF \21mux_2\: COMPONENT IS true;

COMPONENT \21mux_4\
	PORT(S : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 A : IN STD_LOGIC;
		 Y : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \21mux_4\: COMPONENT IS true;
ATTRIBUTE noopt OF \21mux_4\: COMPONENT IS true;

COMPONENT \21mux_5\
	PORT(S : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 A : IN STD_LOGIC;
		 Y : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \21mux_5\: COMPONENT IS true;
ATTRIBUTE noopt OF \21mux_5\: COMPONENT IS true;

COMPONENT \21mux_9\
	PORT(S : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 A : IN STD_LOGIC;
		 Y : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \21mux_9\: COMPONENT IS true;
ATTRIBUTE noopt OF \21mux_9\: COMPONENT IS true;

COMPONENT mux41_0
	PORT(S0 : IN STD_LOGIC;
		 D2 : IN STD_LOGIC;
		 S1 : IN STD_LOGIC;
		 D3 : IN STD_LOGIC;
		 D0 : IN STD_LOGIC;
		 INH : IN STD_LOGIC;
		 D1 : IN STD_LOGIC;
		 Q : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF mux41_0: COMPONENT IS true;
ATTRIBUTE noopt OF mux41_0: COMPONENT IS true;

COMPONENT mux41_1
	PORT(S0 : IN STD_LOGIC;
		 D2 : IN STD_LOGIC;
		 S1 : IN STD_LOGIC;
		 D3 : IN STD_LOGIC;
		 D0 : IN STD_LOGIC;
		 INH : IN STD_LOGIC;
		 D1 : IN STD_LOGIC;
		 Q : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF mux41_1: COMPONENT IS true;
ATTRIBUTE noopt OF mux41_1: COMPONENT IS true;

COMPONENT mux41_14
	PORT(S0 : IN STD_LOGIC;
		 D2 : IN STD_LOGIC;
		 S1 : IN STD_LOGIC;
		 D3 : IN STD_LOGIC;
		 D0 : IN STD_LOGIC;
		 INH : IN STD_LOGIC;
		 D1 : IN STD_LOGIC;
		 Q : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF mux41_14: COMPONENT IS true;
ATTRIBUTE noopt OF mux41_14: COMPONENT IS true;

COMPONENT mux41_15
	PORT(S0 : IN STD_LOGIC;
		 D2 : IN STD_LOGIC;
		 S1 : IN STD_LOGIC;
		 D3 : IN STD_LOGIC;
		 D0 : IN STD_LOGIC;
		 INH : IN STD_LOGIC;
		 D1 : IN STD_LOGIC;
		 Q : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF mux41_15: COMPONENT IS true;
ATTRIBUTE noopt OF mux41_15: COMPONENT IS true;

COMPONENT mux41_3
	PORT(S0 : IN STD_LOGIC;
		 D2 : IN STD_LOGIC;
		 S1 : IN STD_LOGIC;
		 D3 : IN STD_LOGIC;
		 D0 : IN STD_LOGIC;
		 INH : IN STD_LOGIC;
		 D1 : IN STD_LOGIC;
		 Q : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF mux41_3: COMPONENT IS true;
ATTRIBUTE noopt OF mux41_3: COMPONENT IS true;

COMPONENT mux41_6
	PORT(S0 : IN STD_LOGIC;
		 D2 : IN STD_LOGIC;
		 S1 : IN STD_LOGIC;
		 D3 : IN STD_LOGIC;
		 D0 : IN STD_LOGIC;
		 INH : IN STD_LOGIC;
		 D1 : IN STD_LOGIC;
		 Q : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF mux41_6: COMPONENT IS true;
ATTRIBUTE noopt OF mux41_6: COMPONENT IS true;

COMPONENT mux41_7
	PORT(S0 : IN STD_LOGIC;
		 D2 : IN STD_LOGIC;
		 S1 : IN STD_LOGIC;
		 D3 : IN STD_LOGIC;
		 D0 : IN STD_LOGIC;
		 INH : IN STD_LOGIC;
		 D1 : IN STD_LOGIC;
		 Q : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF mux41_7: COMPONENT IS true;
ATTRIBUTE noopt OF mux41_7: COMPONENT IS true;

COMPONENT mux41_8
	PORT(S0 : IN STD_LOGIC;
		 D2 : IN STD_LOGIC;
		 S1 : IN STD_LOGIC;
		 D3 : IN STD_LOGIC;
		 D0 : IN STD_LOGIC;
		 INH : IN STD_LOGIC;
		 D1 : IN STD_LOGIC;
		 Q : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF mux41_8: COMPONENT IS true;
ATTRIBUTE noopt OF mux41_8: COMPONENT IS true;

COMPONENT sumador
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 CIN : IN STD_LOGIC;
		 COUT : OUT STD_LOGIC;
		 S : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT sietesegmentos
	PORT(A0 : IN STD_LOGIC;
		 B0 : IN STD_LOGIC;
		 C0 : IN STD_LOGIC;
		 D0 : IN STD_LOGIC;
		 a : OUT STD_LOGIC;
		 b : OUT STD_LOGIC;
		 c : OUT STD_LOGIC;
		 d : OUT STD_LOGIC;
		 e : OUT STD_LOGIC;
		 f : OUT STD_LOGIC;
		 g : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_92 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_93 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_94 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_95 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_96 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_97 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_98 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_99 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_100 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_71 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_72 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_73 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_74 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_75 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_76 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_77 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_78 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_79 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_80 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_81 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_82 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_83 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_84 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_101 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_102 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_89 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_90 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_0 <= '0';
SYNTHESIZED_WIRE_93 <= '1';
SYNTHESIZED_WIRE_5 <= '0';
SYNTHESIZED_WIRE_6 <= '1';
SYNTHESIZED_WIRE_10 <= '0';
SYNTHESIZED_WIRE_11 <= '1';
SYNTHESIZED_WIRE_17 <= '0';
SYNTHESIZED_WIRE_95 <= '1';
SYNTHESIZED_WIRE_22 <= '0';
SYNTHESIZED_WIRE_97 <= '1';
SYNTHESIZED_WIRE_27 <= '0';
SYNTHESIZED_WIRE_28 <= '1';
SYNTHESIZED_WIRE_44 <= '0';
SYNTHESIZED_WIRE_51 <= '0';
SYNTHESIZED_WIRE_53 <= '1';
SYNTHESIZED_WIRE_84 <= '0';
SYNTHESIZED_WIRE_102 <= '1';
SYNTHESIZED_WIRE_89 <= '0';
SYNTHESIZED_WIRE_90 <= '1';



b2v_inst : mux41_0
PORT MAP(S0 => A0,
		 D2 => SYNTHESIZED_WIRE_0,
		 S1 => S0,
		 D3 => SYNTHESIZED_WIRE_92,
		 D0 => SYNTHESIZED_WIRE_93,
		 INH => SYNTHESIZED_WIRE_93,
		 D1 => SYNTHESIZED_WIRE_92,
		 Q => SYNTHESIZED_WIRE_16);


b2v_inst1 : mux41_1
PORT MAP(S0 => A0,
		 D2 => SYNTHESIZED_WIRE_5,
		 S1 => S0,
		 D3 => B0,
		 D0 => B0,
		 INH => SYNTHESIZED_WIRE_6,
		 D1 => SYNTHESIZED_WIRE_92,
		 Q => SYNTHESIZED_WIRE_15);


b2v_inst10 : 21mux_2
PORT MAP(S => S1,
		 B => SYNTHESIZED_WIRE_8,
		 A => SYNTHESIZED_WIRE_9,
		 Y => F2);






SYNTHESIZED_WIRE_101 <= NOT(B2);



b2v_inst16 : mux41_3
PORT MAP(S0 => A1,
		 D2 => SYNTHESIZED_WIRE_10,
		 S1 => S0,
		 D3 => B1,
		 D0 => B1,
		 INH => SYNTHESIZED_WIRE_11,
		 D1 => SYNTHESIZED_WIRE_94,
		 Q => SYNTHESIZED_WIRE_13);


b2v_inst17 : 21mux_4
PORT MAP(S => S1,
		 B => SYNTHESIZED_WIRE_13,
		 A => SYNTHESIZED_WIRE_14,
		 Y => F1);




b2v_inst2 : 21mux_5
PORT MAP(S => S1,
		 B => SYNTHESIZED_WIRE_15,
		 A => SYNTHESIZED_WIRE_16,
		 Y => F0);


b2v_inst20 : mux41_6
PORT MAP(S0 => A1,
		 D2 => SYNTHESIZED_WIRE_17,
		 S1 => S0,
		 D3 => SYNTHESIZED_WIRE_94,
		 D0 => SYNTHESIZED_WIRE_95,
		 INH => SYNTHESIZED_WIRE_95,
		 D1 => SYNTHESIZED_WIRE_94,
		 Q => SYNTHESIZED_WIRE_14);




SYNTHESIZED_WIRE_94 <= NOT(B1);



b2v_inst24 : mux41_7
PORT MAP(S0 => A3,
		 D2 => SYNTHESIZED_WIRE_22,
		 S1 => S0,
		 D3 => SYNTHESIZED_WIRE_96,
		 D0 => SYNTHESIZED_WIRE_97,
		 INH => SYNTHESIZED_WIRE_97,
		 D1 => SYNTHESIZED_WIRE_96,
		 Q => SYNTHESIZED_WIRE_31);


b2v_inst25 : mux41_8
PORT MAP(S0 => A3,
		 D2 => SYNTHESIZED_WIRE_27,
		 S1 => S0,
		 D3 => B3,
		 D0 => B3,
		 INH => SYNTHESIZED_WIRE_28,
		 D1 => SYNTHESIZED_WIRE_96,
		 Q => SYNTHESIZED_WIRE_30);


b2v_inst26 : 21mux_9
PORT MAP(S => S1,
		 B => SYNTHESIZED_WIRE_30,
		 A => SYNTHESIZED_WIRE_31,
		 Y => F3);







SYNTHESIZED_WIRE_96 <= NOT(B3);



SYNTHESIZED_WIRE_57 <= B1 XOR SYNTHESIZED_WIRE_98;


SYNTHESIZED_WIRE_60 <= B2 XOR SYNTHESIZED_WIRE_98;


SYNTHESIZED_WIRE_66 <= B3 XOR SYNTHESIZED_WIRE_98;


SYNTHESIZED_WIRE_98 <= S0 XOR S1;


b2v_inst36 : 21mux_10
PORT MAP(S => SYNTHESIZED_WIRE_99,
		 B => SYNTHESIZED_WIRE_100,
		 A => A0,
		 Y => SYNTHESIZED_WIRE_37);


SYNTHESIZED_WIRE_100 <= NOT(S0);



SYNTHESIZED_WIRE_99 <= NOT(S1);



SYNTHESIZED_WIRE_63 <= SYNTHESIZED_WIRE_37 XOR SYNTHESIZED_WIRE_100;



b2v_inst40 : 21mux_11
PORT MAP(S => SYNTHESIZED_WIRE_99,
		 B => SYNTHESIZED_WIRE_100,
		 A => A1,
		 Y => SYNTHESIZED_WIRE_45);


b2v_inst41 : 21mux_12
PORT MAP(S => SYNTHESIZED_WIRE_99,
		 B => SYNTHESIZED_WIRE_100,
		 A => A2,
		 Y => SYNTHESIZED_WIRE_47);


b2v_inst42 : 21mux_13
PORT MAP(S => SYNTHESIZED_WIRE_99,
		 B => SYNTHESIZED_WIRE_44,
		 A => A3,
		 Y => SYNTHESIZED_WIRE_49);


SYNTHESIZED_WIRE_56 <= SYNTHESIZED_WIRE_45 XOR SYNTHESIZED_WIRE_100;


SYNTHESIZED_WIRE_59 <= SYNTHESIZED_WIRE_47 XOR SYNTHESIZED_WIRE_100;


SYNTHESIZED_WIRE_65 <= SYNTHESIZED_WIRE_49 XOR SYNTHESIZED_WIRE_100;



SYNTHESIZED_WIRE_69 <= SYNTHESIZED_WIRE_51 XOR S0;


SYNTHESIZED_WIRE_72 <= SYNTHESIZED_WIRE_52 XOR S0;


SYNTHESIZED_WIRE_75 <= S0 XOR S0;



SYNTHESIZED_WIRE_78 <= SYNTHESIZED_WIRE_53 XOR S0;


SYNTHESIZED_WIRE_52 <= SYNTHESIZED_WIRE_54 AND SYNTHESIZED_WIRE_55;


SYNTHESIZED_WIRE_54 <= NOT(S1);



SYNTHESIZED_WIRE_55 <= NOT(S0);





b2v_inst56 : sumador
PORT MAP(A => SYNTHESIZED_WIRE_56,
		 B => SYNTHESIZED_WIRE_57,
		 CIN => SYNTHESIZED_WIRE_58,
		 COUT => SYNTHESIZED_WIRE_61,
		 S => SYNTHESIZED_WIRE_71);


b2v_inst57 : sumador
PORT MAP(A => SYNTHESIZED_WIRE_59,
		 B => SYNTHESIZED_WIRE_60,
		 CIN => SYNTHESIZED_WIRE_61,
		 COUT => SYNTHESIZED_WIRE_67,
		 S => SYNTHESIZED_WIRE_74);


SYNTHESIZED_WIRE_64 <= B0 XOR SYNTHESIZED_WIRE_98;


b2v_inst59 : sumador
PORT MAP(A => SYNTHESIZED_WIRE_63,
		 B => SYNTHESIZED_WIRE_64,
		 CIN => cin,
		 COUT => SYNTHESIZED_WIRE_58,
		 S => SYNTHESIZED_WIRE_68);


SYNTHESIZED_WIRE_92 <= NOT(B0);



b2v_inst60 : sumador
PORT MAP(A => SYNTHESIZED_WIRE_65,
		 B => SYNTHESIZED_WIRE_66,
		 CIN => SYNTHESIZED_WIRE_67,
		 COUT => SYNTHESIZED_WIRE_70,
		 S => SYNTHESIZED_WIRE_77);


b2v_inst61 : sumador
PORT MAP(A => SYNTHESIZED_WIRE_68,
		 B => SYNTHESIZED_WIRE_69,
		 CIN => SYNTHESIZED_WIRE_70,
		 COUT => SYNTHESIZED_WIRE_73,
		 S => SYNTHESIZED_WIRE_80);


b2v_inst62 : sumador
PORT MAP(A => SYNTHESIZED_WIRE_71,
		 B => SYNTHESIZED_WIRE_72,
		 CIN => SYNTHESIZED_WIRE_73,
		 COUT => SYNTHESIZED_WIRE_76,
		 S => SYNTHESIZED_WIRE_81);


b2v_inst63 : sumador
PORT MAP(A => SYNTHESIZED_WIRE_74,
		 B => SYNTHESIZED_WIRE_75,
		 CIN => SYNTHESIZED_WIRE_76,
		 COUT => SYNTHESIZED_WIRE_79,
		 S => SYNTHESIZED_WIRE_82);


b2v_inst64 : sumador
PORT MAP(A => SYNTHESIZED_WIRE_77,
		 B => SYNTHESIZED_WIRE_78,
		 CIN => SYNTHESIZED_WIRE_79,
		 COUT => C0,
		 S => SYNTHESIZED_WIRE_83);


b2v_inst65 : sietesegmentos
PORT MAP(A0 => SYNTHESIZED_WIRE_80,
		 B0 => SYNTHESIZED_WIRE_81,
		 C0 => SYNTHESIZED_WIRE_82,
		 D0 => SYNTHESIZED_WIRE_83,
		 a => a,
		 b => b,
		 c => c,
		 d => d,
		 e => e,
		 f => f,
		 g => g);



b2v_inst8 : mux41_14
PORT MAP(S0 => A2,
		 D2 => SYNTHESIZED_WIRE_84,
		 S1 => S0,
		 D3 => SYNTHESIZED_WIRE_101,
		 D0 => SYNTHESIZED_WIRE_102,
		 INH => SYNTHESIZED_WIRE_102,
		 D1 => SYNTHESIZED_WIRE_101,
		 Q => SYNTHESIZED_WIRE_9);


b2v_inst9 : mux41_15
PORT MAP(S0 => A2,
		 D2 => SYNTHESIZED_WIRE_89,
		 S1 => S0,
		 D3 => B2,
		 D0 => B2,
		 INH => SYNTHESIZED_WIRE_90,
		 D1 => SYNTHESIZED_WIRE_101,
		 Q => SYNTHESIZED_WIRE_8);


END bdf_type;